module arbiter();
endmodule